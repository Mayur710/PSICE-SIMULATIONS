*Active High pass filter 
X1 4 3 5 6 7 UA741
Vs 1 0 AC 1
R1 1 2 10k 
R2 7 3 10k
Vp 5 0 DC 5
Vn 6 0 DC -5
C1 2 3 0.01u
V4 4 0 DC 0
.lib nom.lib
.AC Dec 20 1 100k
.probe 
.end