*Astable Multivibrator 
X1 2 1 4 5 3 UA741
C1 1 0 0.1u
R1 2 0 10k
R2 2 3 10K
R 1 3 4.55k
Vp 4 0 DC 10 
Vn 5 0 DC -10
.lib nom.lib 
.tran 1u 4m 0 1u
.probe 
.end