*bjt current mirror
V1 3 0 DC 5V         ; Power Supply (5V)
I1 3 1 DC 100m       ; Reference Current Source (100mA)
R1 3 4 50            ; Resistor in series with the collector of Q1
Q1 4 2 0 npn_transistor1  ; Reference Transistor (Q1), Emitter grounded
Q2 1 2 0 npn_transistor2  ; Mirror Transistor (Q2), Emitter grounded
.model npn_transistor1 npn (Is=1.8104e-15 Bf=100)
.model npn_transistor2 npn (Is=1.8104e-15 Bf=100)

.tran 1m 100m 10m 10m
.probe
.end