*CE amplifier frequency response 
Vs 1 0 AC 1 SIN(0 1m 1k)
Vcc 5 0 DC 12
R1 2 0 10k
R2 5 2 100k
R3 5 3 20k     ;R3 = Rc
R4 4 0 1k      ;R4 = Re
R5 6 0 100k    ;R5 = Rload
C1 1 2 1u
C2 3 6 1u
C3 4 0 20u
Q1 3 2 4 Q12N3904
.model Q12N3904 NPN (IS=6.734E-15 BF=100.0 NF=1.0 VAF=100.0 IKF=0.3 ISE=3.8E-12 NE=1.5 BR=3.0 NR=1.0 VAR=100.0 RE=0.0 RC=0.1 
+CJE=4.5E-12 CJC=5.0E-12 TF=1.0E-10 TR=5.0E-9)
.AC OCT 10 1 1Gig
.op
.probe
.end