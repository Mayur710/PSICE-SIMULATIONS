*Passive All pass filter
V1 1 0 AC 1
R1 1 2 10k
R2 2 0 10k
R3 1 3 10k
C1 3 0 0.1u

.ac dec 20 10 1meg
.probe
.end