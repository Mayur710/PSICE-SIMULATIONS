*Current Mirror using mosfet
V1 5 0 DC 12 
V2 4 0 DC 12
R1 5 3 120
R2 4 1 120
M1 1 1 0 0 nmosfet
M2 3 1 0 0 nmosfet
.model nmosfet NMOS (PHI=0.7 TOX=9.5E-09 XJ=0.2U TPG=1
+VTO=0.7 DELTA=8.8E-01 LD=5E-08 KP=1.56E-04
+U0=420 THETA=2.3E-01 RSH=2.0E+00 GAMMA=0.62
+NSUB=1.40E+17 NFS=7.20E+11 VMAX=1.8E+05 ETA=2.125E-02
+KAPPA=1E-01 CGDO=3.0E-10 CGSO=3.0E-10
+CGBO=4.5E-10 CJ=5.50E-04 MJ=0.6 CJSW=3E-10
+MJSW=0.35 PB=1.1)
.tran 1m 100m 10m 10m
.probe
.end