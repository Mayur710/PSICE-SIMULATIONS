*Inverting Opamp voltage gain
Vin 1 0 SIN(0 1 1k)
V3 3 0 DC 0
R1 1 2 10k
R2 2 6 20k
Vp 4 0 DC 5
Vn 5 0 DC -5
X1 3 2 4 5 6 UA741
.lib nom.lib
.tran 0.01m 4m 0 0.01m
.probe
.end