*Differential Amplifier mosfet
V1 1 0 SIN(0 1m 1k)
M1 2 1 7 7 nmosfet
M2 4 5 7 7 nmosfet
R1 6 2 5k
R2 6 4 5k
I1 7 8 500u
V2 0 8 3.3
V3 6 0 3.3
V4 5 0 SIN(0 1m 1k 0 0 180)
.model nmosfet NMOS (LEVEL=3 L=2e-06 W=0.5 KP=2e-05 RS=0.01 
+ RD=0.01 VTO=3 RDS=1000000 TOX=2e-06 CGSO=4e-11 CGDO=1e-11
+ CBD=1e-09 MJ=0.5 PB=0.8 FC=0.5 RG=5 IS=1e-14 N=1 RB=0.001 PHI=0.6
+ GAMMA=0 DELTA=0 ETA=0 THETA=0 KAPPA=0 VMAX=0� XJ=0� UO=600)
.tran 1m 5m 0 1m 
.probe
.end

*plot v2-v4 for differential output 