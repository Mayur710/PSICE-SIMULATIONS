*Differential Amplifier using BJT
V1 1 0 SIN(0 10m 1k)
V2 7 0 SIN(0 10m 1k 0 0 180)
V3 6 0 DC 12
V4 0 8 DC 12
R1 6 2 10k
R2 6 5 10k
R3 3 8 20k
Q1 2 1 3 npn_transistor1
Q2 5 7 3 npn_transistor2
.model npn_transistor1 npn (Is=1.8104e-15 Bf=100)
.model npn_transistor2 npn (Is=1.8104e-15 Bf=100)
.tran 1m 10m 1m 1m
.probe
.end
*out put will be differential V2-V5