*Low pass filter using R and L 
V 1 0 AC 1
L 1 2 2m
R1 2 0 10
.AC DEC 20 1 10Meg
.probe
.end