*Weighted summer
V1 1 0 sin(0 2 1k)
V2 2 0 sin(0 1 1k)
Vn 6 0 DC -10
Vp 5 0 DC +10

R1 3 1 10k
R2 3 2 2k
Rf 3 4 10k
*this should give output Vo=-(v1+5v2)=7V 

X1 0 3 5 6 4 uA741

.tran 0.01m 5m 0 0.01m
.lib nom.lib
.probe
.end