*Ideal integrator 
Vin 1 0 PULSE(-5 5 0 0 0 0.5m 1m)
V3 3 0 DC 0
R1 1 2 1k
R2 4 2 10K
R3 4 0 10K
C1 4 2 0.1u
Vp 5 0 DC 10
Vn 6 0 DC -10
X1 0 2 5 6 4 UA741
.lib nom.lib
.tran 0.01m 2m 0.01m
.probe
.end