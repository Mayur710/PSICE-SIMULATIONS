*Active Low pass filter 
X1 4 3 5 6 7 UA741
Vs 1 0 AC 1 
V4 4 0 DC 0
Vn 6 0 DC -5
Vp 5 0 DC 5
R1 1 3 1K
R2 7 3 10k
C1 7 3 0.01u
.lib nom.lib
.AC Dec 20 1 100meg
.probe
.end	