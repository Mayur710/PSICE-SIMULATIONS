*Active differentiator
X1 4 3 5 6 7 UA741
V1 1 0 PULSE(-1 1 0 0 0 100U 200U)
Vp 5 0 DC 15
Vn 6 0 DC -15
R1 1 2 1.6k
R2 4 0 1.5k
R3 3 7 16k
C1 2 3 0.01u
C2 3 7 0.001n
.lib nom.lib
.tran 0.01m 5m 0 0.01m
.probe
.end