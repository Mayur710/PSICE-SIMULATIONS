*Differntial Amplifier 
X1 4 3 5 6 7 UA741
V1 1 0 SIN(0 2 1k)
V2 2 0 SIN(0 5 1k)
Vp 5 0 DC 10
Vn 6 0 DC -10
R1 1 3 2k 
R2 3 7 4k
R3 2 4 2k 
R4 4 0 4k
.lib nom.lib
.tran 0.01m 4m 0 0.01m 
.probe
.end