*Non inverting opamp voltage amplifier 
Vin 1 0 SIN(0 1 1k)
R1 2 0 10K
R2 2 3 10K
Vp 5 0 DC 5
Vn 4 0 DC -5
X1 1 2 5 4 3 UA741
.lib nom.lib 
.tran 0.01m 4m 0 0.01m
.probe
.end