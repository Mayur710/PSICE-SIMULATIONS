*All pass active filter 
X1 3 2 4 5 6 UA741
V1 1 0 AC 1
R1 1 2 10k
R2 1 3 10k
Vp 4 0 DC 5
Vn 5 0 DC -5
R3 2 6 10k
R4 6 0 10k
C1 3 0 0.01u
.lib nom.lib
.ac dec 20 10 1meg
.probe 
.end