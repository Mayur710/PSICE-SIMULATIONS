*passive integrator 
V 1 0 PULSE(0 5 0 10u 10u 1m 2m)
R 1 2 10K
C 2 0 0.01u
.tran 0.01m 20m 0 0.01
.probe
.end